/*MÓDULO RESPONSÁVEL POR TRATAR O RUIDO DO BOTÃO*/
module tratar_botao(
	input botao, 
	input clock, 
	output botao_saida
	);

reg [2:0] estado = 3'b00;
reg debouncer = 1'b0;

always @(posedge clock) begin
	case (estado)
		3'b00: begin
			if(!botao) estado <= estado + 1'b1;
		end
		3'b01: begin
			if(!botao) estado <= estado + 1'b1;
			else estado <= 3'b00;
		end
		3'b10: begin 
			if(!botao) begin
				estado <= estado + 1'b1;
				debouncer <= 1'b1;
			end
			else estado <= 3'b00;
		end
		3'b11: begin
			if(botao) begin
				estado <= 3'b00;
				debouncer <= 1'b0;
			end
		end
	endcase			
end

assign botao_saida = debouncer;
endmodule
